CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 110 10
176 80 1534 813
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100498 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 989 179 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.89883e-315 0
0
2 +V
167 294 256 0 1 3
0 16
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
43529.7 0
0
7 Pulser~
4 195 300 0 10 12
0 18 19 12 12 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
43529.7 1
0
9 CC 7-Seg~
183 1002 238 0 17 19
10 10 9 8 7 6 5 4 20 2
0 1 1 0 0 0 0 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3421 0 0
2
43529.7 2
0
9 2-In AND~
219 684 226 0 3 22
0 3 11 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8157 0 0
2
43529.7 3
0
9 2-In AND~
219 523 224 0 3 22
0 15 14 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43529.7 4
0
6 74112~
219 757 335 0 7 32
0 16 17 12 17 16 21 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
43529.7 5
0
6 74112~
219 610 333 0 7 32
0 16 3 12 22 16 11 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7361 0 0
2
43529.7 6
0
6 74112~
219 441 336 0 7 32
0 16 15 12 15 16 23 14
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4747 0 0
2
43529.7 7
0
6 74112~
219 294 336 0 7 32
0 16 16 12 16 16 24 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
972 0 0
2
43529.7 8
0
6 74LS48
188 893 335 0 14 29
0 13 11 14 15 25 26 4 5 6
7 8 9 10 27
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
43529.7 9
0
37
7 1 0 0 0 0 0 7 11 0 0 2
781 299
861 299
3 1 3 0 0 4224 0 6 5 0 0 4
544 224
652 224
652 217
660 217
7 7 4 0 0 4224 0 11 4 0 0 3
925 299
1017 299
1017 274
8 6 5 0 0 4224 0 11 4 0 0 3
925 308
1011 308
1011 274
9 5 6 0 0 4224 0 11 4 0 0 3
925 317
1005 317
1005 274
10 4 7 0 0 4224 0 11 4 0 0 3
925 326
999 326
999 274
11 3 8 0 0 4224 0 11 4 0 0 3
925 335
993 335
993 274
12 2 9 0 0 4224 0 11 4 0 0 3
925 344
987 344
987 274
13 1 10 0 0 8320 0 11 4 0 0 3
925 353
981 353
981 274
1 9 2 0 0 8320 0 1 4 0 0 3
989 173
1002 173
1002 196
6 0 11 0 0 4096 0 8 0 0 13 2
640 315
641 315
4 0 12 0 0 0 0 3 0 0 25 2
225 300
225 300
0 2 11 0 0 8320 0 0 11 29 0 5
641 297
641 406
837 406
837 308
861 308
0 3 14 0 0 8320 0 0 11 28 0 5
483 300
483 414
847 414
847 317
861 317
0 4 15 0 0 8336 0 0 11 37 0 5
333 300
333 424
856 424
856 326
861 326
0 1 16 0 0 8192 0 0 2 26 0 4
256 300
256 273
294 273
294 265
1 0 16 0 0 0 0 2 0 0 21 2
294 265
294 265
0 0 16 0 0 4096 0 0 0 21 24 2
355 265
355 356
1 1 16 0 0 8192 0 8 7 0 0 4
610 270
610 265
757 265
757 272
1 1 16 0 0 8320 0 9 8 0 0 4
441 273
441 265
610 265
610 270
1 1 16 0 0 0 0 10 9 0 0 4
294 273
294 265
441 265
441 273
5 5 16 0 0 0 0 8 7 0 0 4
610 345
610 356
757 356
757 347
5 5 16 0 0 0 0 9 8 0 0 4
441 348
441 356
610 356
610 345
5 5 16 0 0 0 0 10 9 0 0 4
294 348
294 356
441 356
441 348
3 0 12 0 0 8192 0 3 0 0 34 4
219 291
225 291
225 398
242 398
4 2 16 0 0 0 0 10 10 0 0 4
270 318
256 318
256 300
270 300
2 3 3 0 0 0 0 8 6 0 0 4
586 297
548 297
548 224
544 224
2 7 14 0 0 0 0 6 9 0 0 4
499 233
492 233
492 300
465 300
2 7 11 0 0 0 0 5 8 0 0 4
660 235
652 235
652 297
634 297
2 0 17 0 0 4096 0 7 0 0 31 2
733 299
712 299
3 4 17 0 0 8320 0 5 7 0 0 4
705 226
712 226
712 317
733 317
3 0 12 0 0 0 0 8 0 0 34 3
580 306
554 306
554 399
3 0 12 0 0 0 0 9 0 0 34 3
411 309
397 309
397 399
3 3 12 0 0 12416 0 10 7 0 0 6
264 309
242 309
242 399
702 399
702 308
727 308
1 0 15 0 0 0 0 6 0 0 36 3
499 215
367 215
367 300
4 0 15 0 0 0 0 9 0 0 37 3
417 318
367 318
367 300
7 2 15 0 0 0 0 10 9 0 0 2
318 300
417 300
3
-21 0 0 0 400 0 0 0 0 3 2 1 2
9 DISCOVERY
0 0 0 52
166 93 1081 127
174 100 1072 124
52 FOUR BIT Synchronous Counter Waveform Timing Diagram
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
27 42 116 63
35 48 107 63
9 BSCpE 1-B
-21 0 0 0 700 0 0 0 0 3 2 1 34
14 Century Gothic
0 0 0 23
27 13 312 45
35 20 303 44
23 JAPSON, KITT CYMONNE G.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
